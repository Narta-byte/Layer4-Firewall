library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package my_types_pkg is
    type tree_array is array (natural range <>) of integer;
end package my_types_pkg;
